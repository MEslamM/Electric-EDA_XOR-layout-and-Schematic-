*** SPICE deck for cell XOR_schem{sch} from library XOR
*** Created on Mon May 09, 2022 21:58:38
*** Last revised on Thu May 12, 2022 14:09:31
*** Written on Sun May 22, 2022 20:28:13 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: XOR_schem{sch}
Mnmos@0 net@252 A net@257 gnd NMOS L=0.4U W=1U
Mnmos@1 net@257 B gnd gnd NMOS L=0.4U W=1U
Mnmos@10 net@271 net@252 net@258 gnd NMOS L=0.4U W=1U
Mnmos@11 net@258 A gnd gnd NMOS L=0.4U W=1U
Mnmos@12 net@255 net@252 net@259 gnd NMOS L=0.4U W=1U
Mnmos@13 net@259 B gnd gnd NMOS L=0.4U W=1U
Mnmos@14 Q net@255 net@260 gnd NMOS L=0.4U W=1U
Mnmos@15 net@260 net@271 gnd gnd NMOS L=0.4U W=1U
Mpmos@0 vdd A net@252 vdd PMOS L=0.4U W=2U
Mpmos@1 vdd B net@252 vdd PMOS L=0.4U W=2U
Mpmos@10 vdd net@252 net@271 vdd PMOS L=0.4U W=2U
Mpmos@11 vdd A net@271 vdd PMOS L=0.4U W=2U
Mpmos@12 vdd net@252 net@255 vdd PMOS L=0.4U W=2U
Mpmos@13 vdd B net@255 vdd PMOS L=0.4U W=2U
Mpmos@14 vdd net@255 Q vdd PMOS L=0.4U W=2U
Mpmos@15 vdd net@271 Q vdd PMOS L=0.4U W=2U

* Spice Code nodes in cell cell 'XOR_schem{sch}'
vdd vdd 0 DC 5
va A 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb B 0 DC pwl 10n 0 20n 5 100n 5 110n 0
.tran 200n
.include C:\electric\C5_models.txt
.END
